package beehive_vr_pkg;
    localparam INT_W = 64;
    localparam COUNT_W = 64;

    localparam [31:0]   NONFRAG_MAGIC = 31'h18_03_05_20;

    localparam FRAG_MAGIC_W = 32;
    localparam MSG_LEN_W = 64;

    localparam LOG_W = 512;
    localparam LOG_W_BYTES = LOG_W/8;
    localparam LOG_W_BYTES_W = $clog2(LOG_W_BYTES);
    localparam LOG_DEPTH = 2048;
    localparam LOG_DEPTH_W = $clog2(LOG_DEPTH);
    localparam LOG_HDR_DEPTH = 4096;
    localparam LOG_HDR_DEPTH_W = $clog2(LOG_HDR_DEPTH);

    localparam LOG_STATE_COMMITED = 0;
    localparam LOG_STATE_PREPARED = 1;

    typedef enum logic[7:0] {
        Prepare = 8'd5,
        PrepareOK = 8'd6,
        Commit = 8'd7,
        RequestStateTransfer= 8'd8,
        StateTransfer = 8'd9,
        StartViewChange = 8'd10,
        DoViewChange = 8'd11,
        StartView = 8'd12,
        SetupBeehive = 8'd128
    } msg_type;

    typedef struct packed {
        logic   [FRAG_MAGIC_W-1:0]  frag_num;
        msg_type                    msg_type;
        logic   [MSG_LEN_W-1:0]     msg_len;
    } beehive_hdr;
    localparam BEEHIVE_HDR_W = $bits(beehive_hdr);
    localparam BEEHIVE_HDR_BYTES = BEEHIVE_HDR_W/8;

    typedef struct packed {
        logic   [INT_W-1:0]     view;
        logic   [INT_W-1:0]     opnum;
        logic   [INT_W-1:0]     batchstart;
        logic   [INT_W-1:0]     clean_up_to;
        logic   [COUNT_W-1:0]   req_count;
    } prepare_msg_hdr;
    localparam PREPARE_MSG_HDR_W = $bits(prepare_msg_hdr);
    localparam PREPARE_HDR_BYTES = PREPARE_MSG_HDR_W/8;

    typedef struct packed {
        logic   [INT_W-1:0] view;
        logic   [INT_W-1:0] opnum;
        logic   [INT_W-1:0] rep_index;
        logic   [INT_W-1:0] last_committed;
    } prepare_ok_hdr;
    localparam PREPARE_OK_HDR_W = $bits(prepare_ok_hdr);
    localparam PREPARE_OK_HDR_BYTES = PREPARE_OK_HDR_W/8;

    typedef struct packed {
        logic   [INT_W-1:0]     view;
        logic   [INT_W-1:0]     opnum;
    } commit_msg_hdr;
    localparam COMMIT_MSG_HDR_W = $bits(commit_msg_hdr);

    typedef struct packed {
        logic   [INT_W-1:0]         curr_view;
        logic   [INT_W-1:0]         last_op;
        logic   [INT_W-1:0]         my_replica_index;
        logic   [INT_W-1:0]         first_log_op;
        logic   [LOG_HDR_DEPTH_W:0] hdr_log_head;
        logic   [LOG_HDR_DEPTH_W:0] hdr_log_tail;
        logic   [LOG_DEPTH_W:0]     data_log_head;
        logic   [LOG_DEPTH_W:0]     data_log_tail;
        logic   [INT_W-1:0]         last_commit;
    } vr_state;
    localparam VR_STATE_W = $bits(vr_state);

    typedef struct packed {
        logic   [INT_W-1:0]         view;
        logic   [INT_W-1:0]         op_num;
        logic   [INT_W-1:0]         log_entry_state;
        logic   [INT_W-1:0]         payload_len;
        logic   [LOG_DEPTH_W-1:0]   payload_addr;
        logic   [INT_W-1:0]         req_count;
    } log_entry_hdr;
    localparam LOG_ENTRY_HDR_W = $bits(log_entry_hdr);



endpackage
